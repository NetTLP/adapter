module eth_pcspma_conf (
    output wire [535:0] pcspma_configuration_vector
);
	assign pcspma_configuration_vector = 536'b0;

endmodule

