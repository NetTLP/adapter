module ila_0 (
	input wire clk,
	input wire probe0,
	input wire probe1,
	input wire probe2,
	input wire probe3,
	input wire [1:0] probe4
//	input wire probe5,
//	input wire probe6,
//	input wire probe7,
//	input wire probe8,
//	input wire probe9,
//	input wire probe10,
//	input wire probe11,
//	input wire probe12,
//	input wire probe13
);

wire _unused_ok = &{
	1'b0,
	clk,
	probe0,
	probe1,
	probe2,
	probe3,
	probe4,
//	probe5,
//	probe6,
//	probe7,
//	probe8,
//	probe9,
//	probe10,
//	probe11,
//	probe12,
//	probe13,
	1'b0
};

endmodule

