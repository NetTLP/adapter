module OBUF (
	input  logic I,
	output logic O
);

assign O = I; 

endmodule

