module ila_0 #(
	parameter ILA_PROBE0_WIDTH = 79,
	parameter ILA_PROBE1_WIDTH = 97
)(
	input wire clk,
	input wire [ILA_PROBE0_WIDTH-1:0] probe0,
	input wire [ILA_PROBE1_WIDTH-1:0] probe1
);


endmodule

