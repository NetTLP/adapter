module pcs_pma_conf (
    output wire [535:0] pcs_pma_configuration_vector
);
	assign pcs_pma_configuration_vector = 536'b0;

endmodule

